library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM2 is
port(
      address: in std_logic_vector(3 downto 0);
      output : out std_logic_vector(31 downto 0)
);
end ROM2;

architecture arc_ROM2 of ROM2 is
begin

--         HEX7      HEX6     HEX5     HEX4     HEX3     HEX2     HEX1     HEX0

output <= "0000" & "1110" & "0000" & "1010" & "0011" & "1111" & "0110" & "1001" when address = "0000" else
--          0        E        0        A        3       des      6       9

          "1001" & "0010" & "1111" & "0001" & "1100" & "0101" & "1010" & "1110" when address = "0001" else
--          9        2       des       1        C        5       A       E

          "0101" & "0101" & "1000" & "0111" & "0000" & "1001" & "1110" & "0011" when address = "0010" else
--          5        5        8        7        0        9       E       3

          "1110" & "1101" & "0011" & "1111" & "0100" & "0001" & "1000" & "0100" when address = "0011" else
--          E        D        3       des       4        1       8       4

          "0011" & "1011" & "0100" & "1001" & "1111" & "0111" & "0001" & "0000" when address = "0100" else
--          3        B        4        9       des       7       1       0

          "0110" & "0001" & "1010" & "1100" & "0010" & "1110" & "0101" & "1011" when address = "0101" else
--          6        1        A        C        2        E       5       B

          "1011" & "1000" & "0010" & "0101" & "1010" & "0000" & "1111" & "1100" when address = "0110" else
--          B        8        2        5        A        0      des      C

          "0100" & "1111" & "0111" & "0011" & "1001" & "1010" & "0001" & "0110" when address = "0111" else
--          4       des       7        3        9       A        1       6

          "1100" & "0100" & "1101" & "1000" & "0110" & "0011" & "1011" & "0001" when address = "1000" else
--          C        4        D        8        6        3       B       1

          "0010" & "1010" & "1110" & "0100" & "0001" & "1101" & "1000" & "1111" when address = "1001" else
--          2        A        E        4        1       D       8      des

          "1111" & "0011" & "0001" & "1010" & "0101" & "1000" & "0010" & "0101" when address = "1010" else
--        des        3        1        A        5       8        2       5

          "0001" & "1100" & "0100" & "1110" & "1011" & "0010" & "1100" & "1000" when address = "1011" else
--          1        C        4        E        B        2       C       8

          "0111" & "1001" & "1111" & "0000" & "1100" & "0101" & "0110" & "0010" when address = "1100" else
--          7        9       des       0        C        5       6       2

          "1000" & "0101" & "0011" & "1011" & "1110" & "0001" & "1001" & "0111" when address = "1101" else
--          8        5        3        B        E        1       9       7

          "0100" & "1011" & "0101" & "1100" & "0011" & "1111" & "0000" & "1000" when address = "1110" else
--          4        B        5        C        3       des      0       8

          "1010" & "0000" & "1000" & "0010" & "0111" & "0100" & "1110" & "1101";
--          A        0        8        2        7        4       E       D
end arc_ROM2;