library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM3 is
port(
      address: in std_logic_vector(3 downto 0);
      output : out std_logic_vector(31 downto 0)
);
end ROM3;

architecture arc_ROM3 of ROM3 is
begin

--         HEX7      HEX6     HEX5     HEX4     HEX3     HEX2     HEX1     HEX0

output <= "1110" & "1110" & "0011" & "0001" & "1000" & "0100" & "0101" & "0000" when address = "0000" else
--          E        E        3        1        8        4       5       0

          "0001" & "0011" & "1011" & "0100" & "1110" & "1001" & "1100" & "0111" when address = "0001" else
--          1        3        B        4        E        9       C       7

          "1010" & "0100" & "0001" & "1111" & "0010" & "1100" & "0110" & "1000" when address = "0010" else
--          A        4        1        F        2        C       6       8

          "0111" & "1000" & "0101" & "1011" & "0000" & "0010" & "1111" & "0011" when address = "0011" else
--          7        8        5        B        0        2       F       3

          "0100" & "1010" & "1101" & "0011" & "1001" & "0001" & "1110" & "0101" when address = "0100" else
--          4        A        D        3        9        1       E       5

          "1100" & "0111" & "1001" & "0101" & "0001" & "1010" & "0010" & "1110" when address = "0101" else
--          C        7        9        5        1        A       2       E

          "0010" & "1111" & "0000" & "1100" & "0110" & "0101" & "1000" & "1011" when address = "0110" else
--          2        F        0        C        6        5       8       B

          "1001" & "0000" & "1110" & "0010" & "0101" & "1111" & "0011" & "1100" when address = "0111" else
--          9        0        E        2        5       F       3       C

          "0110" & "1011" & "0010" & "1000" & "1111" & "1101" & "0001" & "0100" when address = "1000" else
--          6        B        2        8        F       D       1       4

          "0100" & "0010" & "0111" & "1100" & "1011" & "1001" & "0001" & "1110" when address = "1001" else
--          4        2        7        C        B       9       1       E

          "1111" & "0010" & "1001" & "0110" & "0100" & "1011" & "0000" & "0011" when address = "1010" else
--          F        2        9        6        4       B       0       3

          "0000" & "1001" & "1110" & "0101" & "1011" & "0011" & "1100" & "0101" when address = "1011" else
--          0        9        E        5        B       3       C       5

          "1011" & "0101" & "1100" & "1111" & "0010" & "0001" & "0110" & "1000" when address = "1100" else
--          B        5        C        F        2       1       6       8

          "0011" & "0110" & "1010" & "1001" & "0001" & "1110" & "0100" & "1011" when address = "1101" else
--          3        6        A        9        1       E       4       B

          "1000" & "1111" & "0100" & "0010" & "0111" & "1010" & "1101" & "0001" when address = "1110" else
--          8        F        4        2        7       A       D       1

          "0100" & "0010" & "0111" & "1100" & "1011" & "1001" & "0001" & "1110";
--          4        2        7        C        B       9       1       E

end arc_ROM3;